`default_nettype none
module genesys_systolic_wrapper #(
  parameter integer C_S_AXI_CONTROL_ADDR_WIDTH    = 12 ,
  parameter integer C_S_AXI_CONTROL_DATA_WIDTH    = 32 ,
  parameter integer C_M00_IMEM_AXI_ADDR_WIDTH     = 64 ,
  parameter integer C_M00_IMEM_AXI_DATA_WIDTH     = 512,
  parameter integer C_M01_PARAMBUF_AXI_ADDR_WIDTH = 64 ,
  parameter integer C_M01_PARAMBUF_AXI_DATA_WIDTH = 512,
  parameter integer C_M02_IBUF_AXI_ADDR_WIDTH     = 64 ,
  parameter integer C_M02_IBUF_AXI_DATA_WIDTH     = 512,
  parameter integer C_M03_OBUF_AXI_ADDR_WIDTH     = 64 ,
  parameter integer C_M03_OBUF_AXI_DATA_WIDTH     = 512
)
(
  input  wire                                       ap_clk                  ,
  input  wire                                       ap_rst_n                ,
  // AXI4 master interface m00_imem_axi
  output wire                                       m00_imem_axi_awvalid    ,
  input  wire                                       m00_imem_axi_awready    ,
  output wire [C_M00_IMEM_AXI_ADDR_WIDTH-1:0]       m00_imem_axi_awaddr     ,
  output wire [8-1:0]                               m00_imem_axi_awlen      ,
  output wire                                       m00_imem_axi_wvalid     ,
  input  wire                                       m00_imem_axi_wready     ,
  output wire [C_M00_IMEM_AXI_DATA_WIDTH-1:0]       m00_imem_axi_wdata      ,
  output wire [C_M00_IMEM_AXI_DATA_WIDTH/8-1:0]     m00_imem_axi_wstrb      ,
  output wire                                       m00_imem_axi_wlast      ,
  input  wire                                       m00_imem_axi_bvalid     ,
  output wire                                       m00_imem_axi_bready     ,
  output wire                                       m00_imem_axi_arvalid    ,
  input  wire                                       m00_imem_axi_arready    ,
  output wire [C_M00_IMEM_AXI_ADDR_WIDTH-1:0]       m00_imem_axi_araddr     ,
  output wire [8-1:0]                               m00_imem_axi_arlen      ,
  input  wire                                       m00_imem_axi_rvalid     ,
  output wire                                       m00_imem_axi_rready     ,
  input  wire [C_M00_IMEM_AXI_DATA_WIDTH-1:0]       m00_imem_axi_rdata      ,
  input  wire                                       m00_imem_axi_rlast      ,
  // AXI4 master interface m01_parambuf_axi
  output wire                                       m01_parambuf_axi_awvalid,
  input  wire                                       m01_parambuf_axi_awready,
  output wire [C_M01_PARAMBUF_AXI_ADDR_WIDTH-1:0]   m01_parambuf_axi_awaddr ,
  output wire [8-1:0]                               m01_parambuf_axi_awlen  ,
  output wire                                       m01_parambuf_axi_wvalid ,
  input  wire                                       m01_parambuf_axi_wready ,
  output wire [C_M01_PARAMBUF_AXI_DATA_WIDTH-1:0]   m01_parambuf_axi_wdata  ,
  output wire [C_M01_PARAMBUF_AXI_DATA_WIDTH/8-1:0] m01_parambuf_axi_wstrb  ,
  output wire                                       m01_parambuf_axi_wlast  ,
  input  wire                                       m01_parambuf_axi_bvalid ,
  output wire                                       m01_parambuf_axi_bready ,
  output wire                                       m01_parambuf_axi_arvalid,
  input  wire                                       m01_parambuf_axi_arready,
  output wire [C_M01_PARAMBUF_AXI_ADDR_WIDTH-1:0]   m01_parambuf_axi_araddr ,
  output wire [8-1:0]                               m01_parambuf_axi_arlen  ,
  input  wire                                       m01_parambuf_axi_rvalid ,
  output wire                                       m01_parambuf_axi_rready ,
  input  wire [C_M01_PARAMBUF_AXI_DATA_WIDTH-1:0]   m01_parambuf_axi_rdata  ,
  input  wire                                       m01_parambuf_axi_rlast  ,
  // AXI4 master interface m02_ibuf_axi
  output wire                                       m02_ibuf_axi_awvalid    ,
  input  wire                                       m02_ibuf_axi_awready    ,
  output wire [C_M02_IBUF_AXI_ADDR_WIDTH-1:0]       m02_ibuf_axi_awaddr     ,
  output wire [8-1:0]                               m02_ibuf_axi_awlen      ,
  output wire                                       m02_ibuf_axi_wvalid     ,
  input  wire                                       m02_ibuf_axi_wready     ,
  output wire [C_M02_IBUF_AXI_DATA_WIDTH-1:0]       m02_ibuf_axi_wdata      ,
  output wire [C_M02_IBUF_AXI_DATA_WIDTH/8-1:0]     m02_ibuf_axi_wstrb      ,
  output wire                                       m02_ibuf_axi_wlast      ,
  input  wire                                       m02_ibuf_axi_bvalid     ,
  output wire                                       m02_ibuf_axi_bready     ,
  output wire                                       m02_ibuf_axi_arvalid    ,
  input  wire                                       m02_ibuf_axi_arready    ,
  output wire [C_M02_IBUF_AXI_ADDR_WIDTH-1:0]       m02_ibuf_axi_araddr     ,
  output wire [8-1:0]                               m02_ibuf_axi_arlen      ,
  input  wire                                       m02_ibuf_axi_rvalid     ,
  output wire                                       m02_ibuf_axi_rready     ,
  input  wire [C_M02_IBUF_AXI_DATA_WIDTH-1:0]       m02_ibuf_axi_rdata      ,
  input  wire                                       m02_ibuf_axi_rlast      ,
  // AXI4 master interface m03_obuf_axi
  output wire                                       m03_obuf_axi_awvalid    ,
  input  wire                                       m03_obuf_axi_awready    ,
  output wire [C_M03_OBUF_AXI_ADDR_WIDTH-1:0]       m03_obuf_axi_awaddr     ,
  output wire [8-1:0]                               m03_obuf_axi_awlen      ,
  output wire                                       m03_obuf_axi_wvalid     ,
  input  wire                                       m03_obuf_axi_wready     ,
  output wire [C_M03_OBUF_AXI_DATA_WIDTH-1:0]       m03_obuf_axi_wdata      ,
  output wire [C_M03_OBUF_AXI_DATA_WIDTH/8-1:0]     m03_obuf_axi_wstrb      ,
  output wire                                       m03_obuf_axi_wlast      ,
  input  wire                                       m03_obuf_axi_bvalid     ,
  output wire                                       m03_obuf_axi_bready     ,
  output wire                                       m03_obuf_axi_arvalid    ,
  input  wire                                       m03_obuf_axi_arready    ,
  output wire [C_M03_OBUF_AXI_ADDR_WIDTH-1:0]       m03_obuf_axi_araddr     ,
  output wire [8-1:0]                               m03_obuf_axi_arlen      ,
  input  wire                                       m03_obuf_axi_rvalid     ,
  output wire                                       m03_obuf_axi_rready     ,
  input  wire [C_M03_OBUF_AXI_DATA_WIDTH-1:0]       m03_obuf_axi_rdata      ,
  input  wire                                       m03_obuf_axi_rlast      ,
  // AXI4 master interface m04_simd_axi
  output wire                                       m04_simd_axi_awvalid    ,
  input  wire                                       m04_simd_axi_awready    ,
  output wire [C_M03_OBUF_AXI_ADDR_WIDTH-1:0]       m04_simd_axi_awaddr     ,
  output wire [8-1:0]                               m04_simd_axi_awlen      ,
  output wire                                       m04_simd_axi_wvalid     ,
  input  wire                                       m04_simd_axi_wready     ,
  output wire [C_M03_OBUF_AXI_DATA_WIDTH-1:0]       m04_simd_axi_wdata      ,
  output wire [C_M03_OBUF_AXI_DATA_WIDTH/8-1:0]     m04_simd_axi_wstrb      ,
  output wire                                       m04_simd_axi_wlast      ,
  input  wire                                       m04_simd_axi_bvalid     ,
  output wire                                       m04_simd_axi_bready     ,
  output wire                                       m04_simd_axi_arvalid    ,
  input  wire                                       m04_simd_axi_arready    ,
  output wire [C_M03_OBUF_AXI_ADDR_WIDTH-1:0]       m04_simd_axi_araddr     ,
  output wire [8-1:0]                               m04_simd_axi_arlen      ,
  input  wire                                       m04_simd_axi_rvalid     ,
  output wire                                       m04_simd_axi_rready     ,
  input  wire [C_M03_OBUF_AXI_DATA_WIDTH-1:0]       m04_simd_axi_rdata      ,
  input  wire                                       m04_simd_axi_rlast      ,
  // Slave Signals
  input  wire                                       s_axi_control_awvalid   ,
  output wire                                       s_axi_control_awready   ,
  input  wire [C_S_AXI_CONTROL_ADDR_WIDTH-1:0]      s_axi_control_awaddr    ,
  input  wire                                       s_axi_control_wvalid    ,
  output wire                                       s_axi_control_wready    ,
  input  wire [C_S_AXI_CONTROL_DATA_WIDTH-1:0]      s_axi_control_wdata     ,
  input  wire [C_S_AXI_CONTROL_DATA_WIDTH/8-1:0]    s_axi_control_wstrb     ,
  input  wire                                       s_axi_control_arvalid   ,
  output wire                                       s_axi_control_arready   ,
  input  wire [C_S_AXI_CONTROL_ADDR_WIDTH-1:0]      s_axi_control_araddr    ,
  output wire                                       s_axi_control_rvalid    ,
  input  wire                                       s_axi_control_rready    ,
  output wire [C_S_AXI_CONTROL_DATA_WIDTH-1:0]      s_axi_control_rdata     ,
  output wire [2-1:0]                               s_axi_control_rresp     ,
  output wire                                       s_axi_control_bvalid    ,
  input  wire                                       s_axi_control_bready    ,
  output wire [2-1:0]                               s_axi_control_bresp     ,
  output wire                                       interrupt               
);

timeunit 1ps;
timeprecision 1ps;

///////////////////////////////////////////////////////////////////////////////
// Parameters
///////////////////////////////////////////////////////////////////////////////

// genesys systolic configuration
`include "config.vh"


///////////////////////////////////////////////////////////////////////////////
// Wires and Variables
///////////////////////////////////////////////////////////////////////////////
(* KEEP = "yes" *)
logic                                areset                         = 1'b0;

///////////////////////////////////////////////////////////////////////////////
// Genesys Accelerator
///////////////////////////////////////////////////////////////////////////////

// Register and invert reset signal.
always @(posedge ap_clk) begin
  areset <= ~ap_rst_n;
end

genesys_top_module #(
    .NUM_TAGS                     (NUM_TAGS               ),      
    .TAG_W                        (TAG_W                  ),  
    .TAG_REUSE_COUNTER_W          (TAG_REUSE_COUNTER_W    ),    
    .ADDR_WIDTH                   (ADDR_WIDTH              ),  
    .ARRAY_N                      (ARRAY_N                ),        
    .ARRAY_M                      (ARRAY_M                ),            
    .DATA_WIDTH                   (DATA_WIDTH             ),                
    .BIAS_WIDTH                   (BIAS_WIDTH             ),                  
    .ACC_WIDTH                    (ACC_WIDTH              ),                
    .IBUF_CAPACITY_BITS           (IBUF_CAPACITY_BITS     ),                            
    .WBUF_CAPACITY_BITS           (WBUF_CAPACITY_BITS     ),                                                                                    
    .OBUF_CAPACITY_BITS           (OBUF_CAPACITY_BITS     ),
    .BBUF_CAPACITY_BITS           (BBUF_CAPACITY_BITS     ),        
    //.IBUF_TAG_ADDR_WIDTH          (IBUF_TAG_ADDR_WIDTH    ),          
    //.OBUF_TAG_ADDR_WIDTH          (OBUF_TAG_ADDR_WIDTH    ),              
    //.WBUF_TAG_ADDR_WIDTH          (WBUF_TAG_ADDR_WIDTH    ),              
    //.BBUF_TAG_ADDR_WIDTH          (BBUF_TAG_ADDR_WIDTH    ),        
    //.IBUF_ADDR_WIDTH              (IBUF_ADDR_WIDTH        ),                                
    //.WBUF_ADDR_WIDTH              (WBUF_ADDR_WIDTH        ),                                
    //.OBUF_ADDR_WIDTH              (OBUF_ADDR_WIDTH        ),                                
    //.BBUF_ADDR_WIDTH              (BBUF_ADDR_WIDTH        ),                                
    //.WBUF_REQ_WIDTH               (WBUF_REQ_WIDTH         ),
    .OBUF_BANK_DEPTH              (OBUF_DEPTH),
    .IBUF_BANK_DEPTH              (IBUF_DEPTH), 
    .WBUF_BANK_DEPTH              (WBUF_DEPTH),
    .BBUF_BANK_DEPTH              (BBUF_DEPTH), 
    .VMEM_ADDR_WIDTH              (VMEM_ADDR_WIDTH),   
    .IMM_ADDR_WIDTH               (IMM_ADDR_WIDTH),
    .SIMD_OPCODE_BITS             (SIMD_OPCODE_BITS), 
    .SIMD_INTERLEAVE              (SIMD_INTERLEAVE),
    .SIMD_FUNCTION_BITS           (SIMD_FUNCTION_BITS), 
    .SIMD_IMEM_ADDR_WIDTH         (SIMD_IMEM_ADDR_WIDTH),                         
    .INST_DATA_WIDTH              (INST_DATA_WIDTH        ),        
    .INST_MEM_CAPACITY_BITS       (INST_MEM_CAPACITY_BITS ),          
    .INST_MEM_ADDR_WIDTH          (INST_MEM_ADDR_WIDTH    ),      
    .BUF_TYPE_W                   (BUF_TYPE_W             ),      
    .IMM_WIDTH                    (IMM_WIDTH              ),        
    .OP_CODE_W                    (OP_CODE_W              ),      
    .OP_SPEC_W                    (OP_SPEC_W              ),      
    .LOOP_ID_W                    (LOOP_ID_W              ),      
    .INST_GROUP_ID_W              (INST_GROUP_ID_W        ),      
    .LOOP_ITER_W                  (LOOP_ITER_W            ),              
    .ADDR_STRIDE_W                (ADDR_STRIDE_W          ),                
    .MEM_REQ_W                    (MEM_REQ_W              ),              
    .GROUP_ENABLED                (GROUP_ENABLED          ),      
    .AXI_ADDR_WIDTH               (AXI_ADDR_WIDTH         ),                
    .AXI_ID_WIDTH                 (AXI_ID_WIDTH           ),      
    .AXI_BURST_WIDTH              (AXI_BURST_WIDTH        ),      
    .INST_MEM_AXI_DATA_WIDTH      (INST_MEM_AXI_DATA_WIDTH),        
    .INST_WSTRB_WIDTH             (INST_WSTRB_WIDTH       ),                                
    .IBUF_AXI_DATA_WIDTH          (IBUF_AXI_DATA_WIDTH    ),        
    .IBUF_WSTRB_WIDTH             (IBUF_WSTRB_WIDTH       ),                            
    .PARAMBUF_AXI_DATA_WIDTH      (PARAMBUF_AXI_DATA_WIDTH),        
    .PARAMBUF_WSTRB_WIDTH         (PARAMBUF_WSTRB_WIDTH   ),                                
    .OBUF_AXI_DATA_WIDTH          (OBUF_AXI_DATA_WIDTH    ),        
    .OBUF_WSTRB_WIDTH             (OBUF_WSTRB_WIDTH       ),                            
    .CTRL_ADDR_WIDTH              (CTRL_ADDR_WIDTH        ),        
    .CTRL_DATA_WIDTH              (CTRL_DATA_WIDTH        ),        
    .CTRL_WSTRB_WIDTH             (CTRL_WSTRB_WIDTH       )                      
) inst_genesys_top_module (

    .clk                       (ap_clk                    ),                          
    .reset                     (areset                    ),                                          
    .pci_cl_ctrl_awvalid       (s_axi_control_awvalid     ),                                          
    .pci_cl_ctrl_awaddr        (s_axi_control_awaddr      ),                                         
    .pci_cl_ctrl_awready       (s_axi_control_awready     ),                                          
    .pci_cl_ctrl_wvalid        (s_axi_control_wvalid      ),                                         
    .pci_cl_ctrl_wdata         (s_axi_control_wdata       ),                                          
    .pci_cl_ctrl_wstrb         (s_axi_control_wstrb       ),                                          
    .pci_cl_ctrl_wready        (s_axi_control_wready      ),                                         
    .pci_cl_ctrl_bvalid        (s_axi_control_bvalid      ),
    .pci_cl_ctrl_bresp         (s_axi_control_bresp       ),                                                                                
    .pci_cl_ctrl_bready        (s_axi_control_bready      ),                                         
    .pci_cl_ctrl_arvalid       (s_axi_control_arvalid     ),                                          
    .pci_cl_ctrl_araddr        (s_axi_control_araddr      ),                                         
    .pci_cl_ctrl_arready       (s_axi_control_arready     ),                                          
    .pci_cl_ctrl_rvalid        (s_axi_control_rvalid      ),
    .pci_cl_ctrl_rresp         (s_axi_control_rresp       ),                                         
    .pci_cl_ctrl_rdata         (s_axi_control_rdata       ),                                                                                  
    .pci_cl_ctrl_rready        (s_axi_control_rready      ),
    .interrupt                 (interrupt                 ),                                                 
    .imem_awaddr               (m00_imem_axi_awaddr       ),                                                  
    .imem_awlen                (m00_imem_axi_awlen        ),                                                                                 
    .imem_awvalid              (m00_imem_axi_awvalid      ),                                           
    .imem_awready              (m00_imem_axi_awready      ),                                            
    .imem_wdata                (m00_imem_axi_wdata        ),                                           
    .imem_wstrb                (m00_imem_axi_wstrb        ),                                           
    .imem_wlast                (m00_imem_axi_wlast        ),                                            
    .imem_wvalid               (m00_imem_axi_wvalid       ),                                             
    .imem_wready               (m00_imem_axi_wready       ),                                                                                      
    .imem_bvalid               (m00_imem_axi_bvalid       ),                                            
    .imem_bready               (m00_imem_axi_bready       ),                                            
    .imem_araddr               (m00_imem_axi_araddr       ),                                           
    .imem_arlen                (m00_imem_axi_arlen        ),                                                                                   
    .imem_arvalid              (m00_imem_axi_arvalid      ),                                                                                     
    .imem_arready              (m00_imem_axi_arready      ),                                            
    .imem_rdata                (m00_imem_axi_rdata        ),                                                                                   
    .imem_rlast                (m00_imem_axi_rlast        ),                                           
    .imem_rvalid               (m00_imem_axi_rvalid       ),                                                                                      
    .imem_rready               (m00_imem_axi_rready       ),                                             
    .parambuf_awaddr           (m01_parambuf_axi_awaddr   ),                                          
    .parambuf_awlen            (m01_parambuf_axi_awlen    ),                                                                                  
    .parambuf_awvalid          (m01_parambuf_axi_awvalid  ),                                         
    .parambuf_awready          (m01_parambuf_axi_awready  ),                                         
    .parambuf_wdata            (m01_parambuf_axi_wdata    ),                                         
    .parambuf_wstrb            (m01_parambuf_axi_wstrb    ),                                         
    .parambuf_wlast            (m01_parambuf_axi_wlast    ),                                         
    .parambuf_wvalid           (m01_parambuf_axi_wvalid   ),                                          
    .parambuf_wready           (m01_parambuf_axi_wready   ),                                                                                  
    .parambuf_bvalid           (m01_parambuf_axi_bvalid   ),                                          
    .parambuf_bready           (m01_parambuf_axi_bready   ),                                          
    .parambuf_araddr           (m01_parambuf_axi_araddr   ),                                                                                   
    .parambuf_arlen            (m01_parambuf_axi_arlen    ),                                                                                  
    .parambuf_arvalid          (m01_parambuf_axi_arvalid  ),                                         
    .parambuf_arready          (m01_parambuf_axi_arready  ),                                         
    .parambuf_rdata            (m01_parambuf_axi_rdata    ),                                                                                                                        
    .parambuf_rlast            (m01_parambuf_axi_rlast    ),                                         
    .parambuf_rvalid           (m01_parambuf_axi_rvalid   ),                                          
    .parambuf_rready           (m01_parambuf_axi_rready   ),                                          
    .ibuf_awaddr               (m02_ibuf_axi_awaddr       ),                                          
    .ibuf_awlen                (m02_ibuf_axi_awlen        ),                                                                                 
    .ibuf_awvalid              (m02_ibuf_axi_awvalid      ),                                         
    .ibuf_awready              (m02_ibuf_axi_awready      ),                                         
    .ibuf_wdata                (m02_ibuf_axi_wdata        ),                                         
    .ibuf_wstrb                (m02_ibuf_axi_wstrb        ),                                         
    .ibuf_wlast                (m02_ibuf_axi_wlast        ),                                         
    .ibuf_wvalid               (m02_ibuf_axi_wvalid       ),                                          
    .ibuf_wready               (m02_ibuf_axi_wready       ),                                                                                  
    .ibuf_bvalid               (m02_ibuf_axi_bvalid       ),                                          
    .ibuf_bready               (m02_ibuf_axi_bready       ),                                          
    .ibuf_araddr               (m02_ibuf_axi_araddr       ),                                          
    .ibuf_arlen                (m02_ibuf_axi_arlen        ),                                                                             
    .ibuf_arvalid              (m02_ibuf_axi_arvalid      ),                                                                        
    .ibuf_arready              (m02_ibuf_axi_arready      ),                                         
    .ibuf_rdata                (m02_ibuf_axi_rdata        ),                                                                                 
    .ibuf_rlast                (m02_ibuf_axi_rlast        ),                                         
    .ibuf_rvalid               (m02_ibuf_axi_rvalid       ),                                                                                  
    .ibuf_rready               (m02_ibuf_axi_rready       ),                                          
    .obuf_awaddr               (m03_obuf_axi_awaddr       ),                                          
    .obuf_awlen                (m03_obuf_axi_awlen        ),                                                                          
    .obuf_awvalid              (m03_obuf_axi_awvalid      ),                                         
    .obuf_awready              (m03_obuf_axi_awready      ),                                         
    .obuf_wdata                (m03_obuf_axi_wdata        ),                                         
    .obuf_wstrb                (m03_obuf_axi_wstrb        ),                                         
    .obuf_wlast                (m03_obuf_axi_wlast        ),                                         
    .obuf_wvalid               (m03_obuf_axi_wvalid       ),                                          
    .obuf_wready               (m03_obuf_axi_wready       ),                                                                                  
    .obuf_bvalid               (m03_obuf_axi_bvalid       ),                                          
    .obuf_bready               (m03_obuf_axi_bready       ),                                          
    .obuf_araddr               (m03_obuf_axi_araddr       ),                                                                                    
    .obuf_arlen                (m03_obuf_axi_arlen        ),                                                                                 
    .obuf_arvalid              (m03_obuf_axi_arvalid      ),                                         
    .obuf_arready              (m03_obuf_axi_arready      ),                                         
    .obuf_rdata                (m03_obuf_axi_rdata        ),                                                                                                                        
    .obuf_rlast                (m03_obuf_axi_rlast        ),                                         
    .obuf_rvalid               (m03_obuf_axi_rvalid       ),                                          
    .obuf_rready               (m03_obuf_axi_rready       ),
    .simd_awaddr               (m04_simd_axi_awaddr       ),                                          
    .simd_awlen                (m04_simd_axi_awlen        ),                                                                          
    .simd_awvalid              (m04_simd_axi_awvalid      ),                                         
    .simd_awready              (m04_simd_axi_awready      ),                                         
    .simd_wdata                (m04_simd_axi_wdata        ),                                         
    .simd_wstrb                (m04_simd_axi_wstrb        ),                                         
    .simd_wlast                (m04_simd_axi_wlast        ),                                         
    .simd_wvalid               (m04_simd_axi_wvalid       ),                                          
    .simd_wready               (m04_simd_axi_wready       ),                                                                                  
    .simd_bvalid               (m04_simd_axi_bvalid       ),                                          
    .simd_bready               (m04_simd_axi_bready       ),                                          
    .simd_araddr               (m04_simd_axi_araddr       ),                                                                                    
    .simd_arlen                (m04_simd_axi_arlen        ),                                                                                 
    .simd_arvalid              (m04_simd_axi_arvalid      ),                                         
    .simd_arready              (m04_simd_axi_arready      ),                                         
    .simd_rdata                (m04_simd_axi_rdata        ),                                                                                                                        
    .simd_rlast                (m04_simd_axi_rlast        ),                                         
    .simd_rvalid               (m04_simd_axi_rvalid       ),                                          
    .simd_rready               (m04_simd_axi_rready       )                          
);

endmodule : genesys_systolic_wrapper
`default_nettype wire
